package Servo_PKG;

	typedef enum {
		SERVO_POS_UP,
		SERVO_POS_DOWN
	} ServoPos_t;

	typedef enum {
		SERVO_DIR_UP,
		SERVO_DIR_DOWN,
		SERVO_DIR_STAY
	} ServoDir_t;

endpackage : Servo_PKG
