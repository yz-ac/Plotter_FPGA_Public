package Position_PKG;

	typedef enum {
		POS_DIR_UP,
		POS_DIR_DOWN,
		POS_DIR_LEFT,
		POS_DIR_RIGHT
	} PosDirection_t;

	typedef enum {
		POS_QUADRANT_1 = 1,
		POS_QUADRANT_2 = 2,
		POS_QUADRANT_3 = 3,
		POS_QUADRANT_4 = 4
	} PosQuadrant_t;

endpackage : Position_PKG
