`ifndef __OP_SVH__
`define __OP_SVH__

`define OP_BITS (64)
`define OP_ARG_BITS (12)
`define OP_CMD_BITS (8)
`define OP_ARG_1_BITS (`OP_ARG_BITS)
`define OP_ARG_2_BITS (`OP_ARG_BITS)
`define OP_ARG_3_BITS (`OP_ARG_BITS)
`define OP_ARG_4_BITS (`OP_ARG_BITS)
`define OP_FLAGS_BITS (8)

`define OP_FLAGS_AXES_CROSS_BIT (0)
`define OP_FLAGS_FULL_CIRCLE_BIT (1)

`endif // __OP_SVH__
