`ifndef __TYPES_SVH__
`define __TYPES_SVH__

`define NIBBLE_BITS (4)
`define BYTE_BITS (8)
`define WORD_BITS (16)
`define DWORD_BITS (32)
`define QWORD_BITS (64)

`endif // __TYPES_SVH__
