`ifndef __POSITION_SVH__
`define __POSITION_SVH__

`include "common/common.svh"

`define POS_X_BITS (`OP_ARG_1_BITS)
`define POS_Y_BITS (`OP_ARG_2_BITS)

`endif // __POSITION_SVH__
