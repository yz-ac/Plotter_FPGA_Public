`ifndef __CLOCKING_SVH__
`define __CLOCKING_SVH__

`include "clocking/mmcm.svh"

`endif // __CLOCKING_SVH__
