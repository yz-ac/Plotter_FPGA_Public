`ifndef __PROCESSOR_SVH__
`define __PROCESSOR_SVH__

`include "../../src/common/common.svh"
`include "../../src/common/opcode.svh"

`define STEPPER_X_BITS (`ARG_BITS)
`define STEPPER_Y_BITS (`ARG_BITS)

`endif // __PROCESSOR_SVH__
