`ifndef __MMCM_SVH__
`define __MMCM_SVH__

`define CLKOUT_MULT_F (9.125)
`define CLKOUT_DIV_F (36.500)

`endif // __MMCM_SVH__
