`include "../common/common.svh"

module LinearOpProcessor #(
	ARG_BITS = `ARG_BITS,
	FLAG_BITS = `FLAG_BITS
)
