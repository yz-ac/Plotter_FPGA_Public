package Char_PKG;

	typedef enum {
		CHAR_G,
		CHAR_NUM,
		CHAR_X,
		CHAR_Y,
		CHAR_I,
		CHAR_J,
		CHAR_WHITESPACE,
		CHAR_DOT,
		CHAR_NEWLINE,
		CHAR_UNKNOWN
	} Char_t;

endpackage : Char_PKG
