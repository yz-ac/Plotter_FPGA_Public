`ifndef __OP_SVH__
`define __OP_SVH__

`define OP_CMD_BITS (8)
`define OP_ARG_1_BITS (12)
`define OP_ARG_2_BITS (12)
`define OP_ARG_3_BITS (12)
`define OP_ARG_4_BITS (12)
`define OP_FLAGS_BITS (8)
`define OP_BITS (64)

`endif // __OP_SVH__
