`ifndef __PERIPHERALS_SVH__
`define __PERIPHERALS_SVH__

`include "peripherals/stepper.svh"
`include "peripherals/servo.svh"

`endif // __PERIPHERALS_SVH__
