`ifndef __SIMULATION_SVH__
`define __SIMULATION_SVH__

`timescale 1ns/1ps
`define CLOCK_PERIOD (20) // ns

`define TEST_OUT_FILE "out/tb_test.txt"

`endif // __SIMULATION_SVH__
