`ifndef __UART_SVH__
`define __UART_SVH__

`include "uart/uart_115200_8.svh"

`endif // __UART_SVH__
