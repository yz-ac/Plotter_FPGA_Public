`ifndef __MOTORS_SVH__
`define __MOTORS_SVH__

`include "motors/stepper.svh"
`include "motors/servo.svh"

`endif // __MOTORS_SVH__
