`ifndef __STEPPER_SVH__
`define __STEPPER_SVH__

`include "common/common.svh"

`ifdef SIM_DEBUG

`define STEPPER_PULSE_NUM_X_FACTOR (2)
`define STEPPER_PULSE_NUM_Y_FACTOR (2)


`define STEPPER_PULSE_NUM_X_BITS (`OP_ARG_1_BITS)
`define STEPPER_PULSE_NUM_Y_BITS (`OP_ARG_2_BITS)
`define STEPPER_PULSE_WIDTH_BITS (`BYTE_BITS)
`define STEPPER_PULSE_WIDTH (5)

`else // SIM_DEBUG

`define STEPPER_PULSE_NUM_X_FACTOR (10)
`define STEPPER_PULSE_NUM_Y_FACTOR (10)

`define STEPPER_PULSE_NUM_X_BITS (`OP_ARG_1_BITS)
`define STEPPER_PULSE_NUM_Y_BITS (`OP_ARG_2_BITS)
`define STEPPER_PULSE_WIDTH_BITS (`DWORD_BITS)
`define STEPPER_PULSE_WIDTH (50_000) // 2ms min pulses (40ns clk)

`endif // SIM_DEBUG

`endif // __STEPPER_SVH__
