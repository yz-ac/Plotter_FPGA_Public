`ifndef __VGA_SVH__
`define __VGA_SVH__

`include "vga/vga_640_480_60.svh"

`endif // __VGA_SVH__
