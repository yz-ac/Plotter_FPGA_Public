`ifndef __PROCESSOR_SVH__
`define __PROCESSOR_SVH__

`include "processor/stepper.svh"
`include "processor/servo.svh"

`endif // __PROCESSOR_SVH__
