`ifndef __COMMON_SVH__
`define __COMMON_SVH__

// Standard sizes
`define NIBBLE_BITS (4)
`define BYTE_BITS (8)
`define WORD_BITS (16)
`define DWORD_BITS (32)
`define QWORD_BITS (64)

// Board constants
`define CLOCK_PERIOD (20) // ns

`endif // __COMMON_SVH__
