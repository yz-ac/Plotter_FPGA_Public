`ifndef __PROCESSOR_SVH__
`define __PROCESSOR_SVH__

`include "processor/position.svh"

`endif // __PROCESSOR_SVH__
