package Servo_P;

	typedef enum {
		SERVO_POS_UP,
		SERVO_POS_DOWN
	} ServoPos_t;

	typedef enum {
		SERVO_MOV_UP,
		SERVO_MOV_CENTER,
		SERVO_MOV_DOWN
	} ServoMov_t;

endpackage : Servo_P
