`ifndef __COMMON_SVH__
`define __COMMON_SVH__

`include "common/types.svh"
`include "common/op.svh"

`endif // __COMMON_SVH__
