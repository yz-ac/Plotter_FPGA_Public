`ifndef __COMMON_SVH__
`define __COMMON_SVH__

`include "common/types.svh"

`endif // __COMMON_SVH__
